// 110652011
module Hazard_Detection(clk, )


endmodule